`include "../core/defines.v"

module timer
(
  input clk,
  input rst_n,
  input [31:0] waddr_i,
  input [31:0] wdata_i,
  output [31:0] rdata_o,
  output [31:0] int_req_o
);



endmodule
